package ft232h_package;
    parameter FT232H_AXIS_ASYNC_FIFO_DEPTH = 64;
    parameter FT232H_AXIS_ASYNC_FIFO_DATA_WIDTH = 8;

    parameter FT232H_BFM_AXIS_FIFO_DEPTH = 2;
endpackage